library verilog;
use verilog.vl_types.all;
entity ex4_vlg_tst is
end ex4_vlg_tst;
