library verilog;
use verilog.vl_types.all;
entity ex2_vlg_tst is
end ex2_vlg_tst;
