library verilog;
use verilog.vl_types.all;
entity ex1_vlg_tst is
end ex1_vlg_tst;
