library verilog;
use verilog.vl_types.all;
entity ex12_vlg_tst is
end ex12_vlg_tst;
