library verilog;
use verilog.vl_types.all;
entity ex13_vlg_tst is
end ex13_vlg_tst;
