library verilog;
use verilog.vl_types.all;
entity ex3_vlg_tst is
end ex3_vlg_tst;
