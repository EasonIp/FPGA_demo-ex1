library verilog;
use verilog.vl_types.all;
entity ex6_vlg_tst is
end ex6_vlg_tst;
